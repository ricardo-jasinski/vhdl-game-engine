library ieee;
use ieee.std_logic_1164.all;
use work.basic_types_pkg.all;
use work.input_types_pkg.all;
use work.graphics_types_pkg.all;
use work.sprites_pkg.all;
use work.game_state_pkg.all;
use work.resource_handles_pkg.all;
use work.resource_data_pkg.all;
use work.resource_data_helper_pkg.all;
use work.npc_pkg.all;
use work.vga_pkg.all;

-- Top-level entity for the "Adventure" game demo using VAGE. On top of this
-- entity, there should be only a very simple wrapper intantiating this entity
-- and connecting its ports to the board used. It should be fairly easy to use
-- this entity in other hardware platforms, without any modifications.
entity space_shooter_demo_top is
    port (
        -- synchronous reset, used by all user logic
        reset: in std_logic;
        -- system clock used for all user logic
        clock_50_Mhz: in std_logic;
        -- VGA clock used by the video renderer; should be approximately
        -- 25.715 MHz (25 MHz is acceptable)
        vga_clock_in: in std_logic;
        -- Same as VGA input clock, must be passed along to the video DAC chip
        vga_clock_out: out std_logic;
        -- VGA blank, low during horizontal or vertical retrace (pixels should be blank)
        vga_blank: out std_logic;
        -- VGA Hsync, low during horizontal synchronism pulse
        vga_n_hsync: out std_logic;
        -- VGA Vsync, low during vertical synchronism pulse
        vga_n_vsync: out std_logic;
        -- Composite sync for the ADV7123; if this feature is not used, should
        -- be tied to '0'
        vga_n_sync: out std_logic;
        -- VGA red channel output
        vga_red: out std_logic_vector(9 downto 0);
        -- VGA green channel output
        vga_green: out std_logic_vector(9 downto 0);
        -- VGA blue channel output
        vga_blue: out std_logic_vector(9 downto 0);
        -- Input toggle switches, active high
        input_switches: in std_logic_vector(1 downto 0);
        -- Input push-button switches, active high
        input_buttons: in std_logic_vector(3 downto 0);
        -- Debug pins for debugging game logic (e.g., connecting to board leds)
        debug_bits: out std_logic_vector(7 downto 0)
    );
end;

architecture rtl of space_shooter_demo_top is

    -- Medium-resolution time base (used for game state updates and
    -- reading the inputs switches)
    signal time_base_50_ms: std_logic;
    -- Maximum value for the game time counter
    constant GAME_TIMER_50_MS_MAX: integer := 1000;
    -- Monotonic game time counter, updated every 50 ms. Can be used by
    -- the game logic (eg., to animate or move sprites)
    signal elapsed_time: integer range 0 to GAME_TIMER_50_MS_MAX;

    -- Video engine output uses custom data type; we'll convert here to std_logic
    signal vga_output_signals: vga_output_signals_type;

    -- Array containing the position of each sprite on the screen; generated by
    -- the game logic module and used as an input by the sprites engine
    signal sprite_positions: point_array_type(GAME_SPRITES'range);

    -- We need to tell the sprites engine which sprites we want to monitor for
    -- collisions. The query array helps us do it neatly.
    constant SPRITES_COLLISION_QUERY: sprite_collision_query_type := make_sprites_collision_query((
        (SORCERER_SPRITE, GHOST_SPRITE),
        (SORCERER_SPRITE, SCORPION_SPRITE),
        (SORCERER_SPRITE, ORYX_11_SPRITE),
        (SORCERER_SPRITE, CHEST_SPRITE)
    ));

    -- Each element is 'true' while the two corresponding sprites are colliding.
    signal sprite_collisions: bool_vector(SPRITES_COLLISION_QUERY'range);

    -- We need to initialize the sprites engine with the game sprites. This
    -- initialization array helps us do it neatly. The helper function will
    -- fetch user-provided data from the GAME_SPRITES array and return an
    -- array of sprites ready to be assigned to sprite engine upon reset.
    constant SPRITES_INITIAL_VALUES: sprites_array_type := make_sprites_initial_values(GAME_SPRITES);

    -- Background image to be used by the video engine; currently, the game
    -- logic is responsible for providing the video engine with background tile
    signal background_bitmap: paletted_bitmap_type(0 to 7, 0 to 7);

    -- Define the Non-Player Characters (NPCs) used in the game. The NPCs have
    -- their positions updated automatically; the user logic is responsible for
    -- reading their positions and assigning them to the corresponding sprites
    constant NPCS: npc_array_type := (
        -- Ghost, moves around the chest in a diamond-shaped path
        make_npc_bouncer(
            initial_position => (144, 64),
            allowed_region => (128, 64, 160, 96),
            initial_speed => (1, 1)
        ),
        -- Scorpion, moves horizontally accross the screen
        make_npc_bouncer(
            initial_position => (0, 128),
            initial_speed => (1, 0)
        ),
        -- Bat, moves horizontally
        make_npc_bouncer(
            initial_position => (160, 160),
            allowed_region => (0, 160, 300, 164),
            initial_speed => (1, 1)
        ),
        -- Oryx, tries to kill the player with its sword
        make_npc_follower(
            initial_position => (300, 220),
            slowdown_factor => 2
        ),
        -- Archer, tries to hide behind the player
        make_npc_follower(
            initial_position => (0, 0),
            slowdown_factor => 1
        ),
        -- Reaper, stays near the player
        make_npc_follower(
            initial_position => (300, 64),
            slowdown_factor => 4
        )
    );

    -- User logic must inform the NPC engine what are the target positions
    -- for the NPCs; some types of AI (e.g., AI_FOLLOWER) use this value to
    -- calculate their next position
    signal npc_target_positions: point_array_type(NPCS'range);
    -- The game engine (NPC engine, actually) calculates the NPC positions
    -- and these values are handed over to the game logic
    signal npc_positions: point_array_type(NPCS'range);

    signal in_buttons: input_buttons_type;
    signal game_state: game_state_type;

begin

    ----------------------------------------------------------------------------
    -- Overall architecture description:
    --   1) Instantiate the game logic
    --   2) Instantiate the NPC engine
    --   3) Instantiate the game engine
    --   4) Select a background bitmap based on the current game state
    --   5) Convert signals between std_logic and custom data types. Internally,
    --      we use custom types for better abstraction; at the interface, we use
    --      std_logic for better portability and easier instantiation
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    -- Section 1) Instantiate the game logic. This entity receives the raw game
    -- data and events, and updates the game state accordingly.

    logic: entity work.game_logic
        port map(
            clock => clock_50_Mhz,
            reset => reset,
            time_base_50_ms => time_base_50_ms,
            npc_positions => npc_positions,
            npc_target_positions => npc_target_positions,
            sprite_collisions => sprite_collisions,
            sprites_positions => sprite_positions,
            input_buttons  => in_buttons,
            game_state => game_state,
            debug_bits => debug_bits
        );

    ----------------------------------------------------------------------------
    -- Section 2) Instantiate the NPC engine. This entity receives low-level
    -- game data, and updates the NPC positions.

    npc: entity work.npcs_engine
        generic map (
            NPC_DEFINITIONS => NPCS
        ) port map (
            clock => clock_50_Mhz,
            reset => reset,
            time_base => time_base_50_ms,
            target_positions => npc_target_positions,
            npc_positions => npc_positions
        );

    ----------------------------------------------------------------------------
    -- Section 3) Instantiate the game engine. While game logic performs
    -- functions that are more related with the game itself, the game engine
    -- performs basic functions such as calculating sprite collisions and
    -- rendering the video output.

    engine: entity work.game_engine
        generic map (
            SPRITES_INITIAL_VALUES => SPRITES_INITIAL_VALUES,
            SPRITES_COLLISION_QUERY => SPRITES_COLLISION_QUERY
        ) port map (
            clock_50MHz => clock_50_Mhz,
            reset => reset,
            sprites_coordinates => sprite_positions,
            sprite_collisions_results => sprite_collisions,
            elapsed_time => elapsed_time,
            time_base_50_ms => time_base_50_ms,
            game_state => game_state,
            background_bitmap => background_bitmap,
            vga_clock_in => vga_clock_in,
            vga_signals => vga_output_signals
        );

    ----------------------------------------------------------------------------
    -- Section 4)
    -- Select a background bitmap based on current game state (currently, this
    -- is the only feedback we provide the player with)

    with game_state select background_bitmap <=
        get_bitmap_from_handle(GAME_OVER_TILE_BITMAP) when GS_GAME_OVER,
        get_bitmap_from_handle(GAME_WON_TILE_BITMAP) when GS_GAME_WON,
        get_bitmap_from_handle(FOREST_TILE_BITMAP) when others;

    ----------------------------------------------------------------------------
    -- Section 5) Convert signals between std_logic and custom data types.
    -- Internally, we use custom types for better abstraction; at the interface,
    -- we use std_logic for better portability and easier instantiation.

    -- Connect each pushbutton to the corresponding game input function
    in_buttons <= (
        up => input_buttons(3),
        down => input_buttons(2),
        left => input_buttons(1),
        right => input_buttons(0)
    );

    -- Connect each VGA output signal to the correspoding VGA pin or port
    vga_clock_out <= vga_output_signals.vga_clock_out;
    vga_blank <= vga_output_signals.blank;
    vga_n_hsync <= vga_output_signals.hsync;
    vga_n_vsync <= vga_output_signals.vsync;
    vga_n_sync <= vga_output_signals.sync;
    vga_red <= vga_output_signals.red;
    vga_green <= vga_output_signals.green;
    vga_blue <= vga_output_signals.blue;

end;