package basic_types_pkg is
    type bool_vector is array (natural range <>) of boolean;
end;