package game_state_pkg is
    type game_state_type is (GS_RESET, GS_PLAY, GS_GAME_OVER, GS_GAME_WON);
end;
