use work.sprites_pkg.all;
use work.graphics_types_pkg.all;
use work.resource_handles_pkg.all;
use work.resource_handles_helper_pkg.all;

package resource_data_pkg is

    -- Here we define all the sprites used in the game
    constant GAME_SPRITES: sprite_init_array_type := (
        (SORCERER_SPRITE, bitmap_handle => SORCERER_BITMAP),
        (AXE_SPRITE,      bitmap_handle => AXE_BITMAP     ),
        (ARCHER_SPRITE,   bitmap_handle => ARCHER_BITMAP  ),
        (CHEST_SPRITE,    bitmap_handle => CHEST_BITMAP   ),
        (GHOST_SPRITE,    bitmap_handle => GHOST_BITMAP   ),
        (SCORPION_SPRITE, bitmap_handle => SCORPION_BITMAP),
        (ORYX_11_SPRITE,  bitmap_handle => ORYX_11_BITMAP ),
        (ORYX_12_SPRITE,  bitmap_handle => ORYX_12_BITMAP ),
        (ORYX_21_SPRITE,  bitmap_handle => ORYX_21_BITMAP ),
        (ORYX_22_SPRITE,  bitmap_handle => ORYX_22_BITMAP ),
        (BAT_SPRITE,      bitmap_handle => BAT_BITMAP     ),
        (REAPER_SPRITE,   bitmap_handle => REAPER_BITMAP  )
    );

    -- Here we define the actual bitmaps for each sprite in the game. This is
    -- the second step to add a new sprite in the game.
    constant GAME_BITMAPS: bitmap_init_array_type := (
        (
            handle => SORCERER_BITMAP,
            bitmap => (
                (23, 23, 24, 24, 23,  0, 20, 20),
                ( 0, 23, 24, 24, 23, 23,  0, 20),
                (23, 23, 57, 34, 57, 34,  0, 61),
                ( 0, 23, 23, 57, 57, 57,  0, 20),
                (23, 23, 24, 24, 24, 23, 23, 57),
                (57, 20, 20, 20, 19, 20,  0, 20),
                ( 0, 23, 23, 23, 23, 23,  0, 20),
                (23, 19, 23, 23, 23, 19,  0, 19)
            )
        ),
        (
            handle => AXE_BITMAP,
            bitmap => (
                ( 0,  0,  0,  0,  0,  0,  0,  0),
                ( 0,  0,  0, 18,  0,  0, 37,  0),
                ( 0,  0,  0,  0, 18, 18,  0,  0),
                ( 0,  0,  0,  0, 18, 18, 18, 19),
                ( 0,  0,  0, 37,  0, 18, 19, 19),
                ( 0,  0, 37,  0,  0, 19, 19,  0),
                ( 0, 37,  0,  0,  0,  0,  0,  0),
                (37,  0,  0,  0,  0,  0,  0,  0)
            )
        ),
        (
            handle => ARCHER_BITMAP,
            bitmap => (
                (29, 29, 30, 30, 29,  0, 25,  0),
                ( 0, 29, 30, 30, 30, 29,  0, 25),
                ( 0, 29, 57, 34, 57, 34,  0, 25),
                ( 0,  3, 57, 57, 57, 57,  0, 25),
                (44, 29, 30, 30, 30, 29, 29, 57),
                (57, 37, 38, 38, 19, 37,  0, 41),
                ( 0, 29, 29, 29, 29, 29,  0, 25),
                ( 0, 37,  0,  0,  0, 37, 38,  0)
            )
        ),
        (
            handle => CHEST_BITMAP,
            bitmap => (
                ( 0,  0,  0,  0,  0,  0,  0,  0),
                ( 0, 38, 38, 38, 38, 38, 38,  0),
                (38,  2,  2,  2,  2, 38,  2, 38),
                (38, 38, 38, 38, 38, 38, 38, 38),
                (38,  1, 46,  1, 22, 38, 22, 38),
                (38, 21, 21,  1, 22, 37, 22, 38),
                (37, 37, 37, 37, 37, 37, 37, 37),
                ( 0,  0,  0,  0,  0,  0,  0,  0)
            )
        ),
        (
            handle => GHOST_BITMAP,
            bitmap => (
                ( 0,  0,  0, 53, 53, 53, 20,  0),
                ( 0,  0, 53, 53, 24, 53, 24,  0),
                ( 0,  0, 53, 53, 53, 53, 53,  0),
                ( 0, 53, 53, 53, 53, 34, 53, 53),
                ( 0,  0, 53, 53, 53, 34, 20,  0),
                (53,  0, 53, 53, 53, 53, 20,  0),
                ( 0, 53, 53, 53, 53, 53, 20,  0),
                ( 0,  0, 53, 53, 53, 20,  0,  0)
            )
        ),
        (
            handle => SCORPION_BITMAP,
            bitmap => (
                ( 0, 18, 18, 18,  0,  0,  0,  0),
                (18,  0,  0, 17, 17,  0,  0,  0),
                (18,  0,  0,  0, 17,  0,  0,  0),
                (18,  0,  0,  0,  0,  0,  0,  0),
                (18, 18,  0,  0,  0,  0,  0,  0),
                (17, 18, 18, 18, 18, 24, 18, 24),
                ( 0, 17, 18, 18, 18, 18, 18, 18),
                (17,  0, 17,  0, 17,  0, 17,  0)
            )
        ),
        (
            handle => ORYX_11_BITMAP,
            bitmap => (
                ( 0, 20,  0,  0, 20,  0,  0,  0),
                (20, 20,  0, 20,  0,  0, 34, 34),
                (20, 20,  0, 20,  0, 34, 17, 17),
                (20, 20,  0,  0, 20, 34, 17, 17),
                (20, 20,  0,  0,  0, 33, 24, 34),
                (20, 20,  0,  0, 34, 33, 33, 34),
                (34, 34,  0, 34, 33, 34, 33, 34),
                (17, 34, 17, 34, 17, 33, 34, 33)
            )
        ),
        (
            handle => ORYX_12_BITMAP,
            bitmap => (
                ( 0,  0,  0, 20,  0,  0,  0,  0),
                (34, 34,  0,  0, 20,  0,  0,  0),
                (33, 33, 34,  0, 20,  0,  0,  0),
                (34, 33, 34, 20,  0,  0,  0,  0),
                (34, 24, 33,  0,  0,  0,  0,  0),
                (34, 33, 33, 34,  0,  0,  0,  0),
                (34, 33, 34, 34, 34, 34, 34, 34),
                (33, 34, 17, 34, 18, 18, 18, 34)
            )
        ),
        (
            handle => ORYX_21_BITMAP,
            bitmap => (
                (17, 34, 17, 34, 33, 17, 17, 34),
                (34, 34,  0,  0, 34, 34, 34, 33),
                (34,  0,  0,  0,  0, 34, 33, 33),
                ( 0,  0,  0,  0, 34, 17, 34, 34),
                ( 0,  0,  0, 34, 17, 34, 34, 17),
                ( 0,  0,  0, 34, 34, 34,  0, 33),
                ( 0,  0,  0, 34, 34, 34,  0,  0),
                ( 0,  0, 34, 34, 34, 34,  0,  0)
            )
        ),
        (
            handle => ORYX_22_BITMAP,
            bitmap => (
                (34, 17, 17, 34, 18, 18, 20, 34),
                (33, 34, 34, 34, 18, 20, 20, 34),
                (33, 33, 34, 34, 18, 18, 20, 34),
                (34, 34, 17, 34, 18, 18, 20, 34),
                (17, 34, 34, 17, 34, 18, 18, 34),
                (33,  0, 34, 34, 34, 34, 34, 34),
                ( 0,  0, 34, 34, 34,  0,  0,  0),
                ( 0,  0, 34, 34, 34, 34,  0,  0)
            )
        ),
        (
            handle => BAT_BITMAP,
            bitmap => (
                ( 0,  0,  0, 17,  0, 17,  0,  0),
                ( 0, 17,  0, 17, 17, 17,  0, 17),
                (17, 17,  0, 46, 17, 46,  0, 17),
                (17, 17, 17, 17, 17, 17, 17, 17),
                (17, 17, 17, 17, 17, 17, 17, 17),
                (17, 17,  0, 17, 17,  0, 17, 17),
                (17,  0,  0, 17,  0,  0,  0, 17),
                ( 0,  0,  0,  0,  0,  0,  0,  0)
            )
        ),
       (    handle => REAPER_BITMAP,
            bitmap => (
                (34, 34, 34, 19, 19, 19, 19, 19),
                ( 0, 34, 19, 33, 33, 33,  0, 38),
                ( 0, 34, 34, 23, 53, 23,  0, 38),
                ( 0, 34, 34, 53, 53, 53,  0, 38),
                (34, 34, 34, 34, 34, 34, 34, 53),
                (53, 34, 34, 34, 34, 34,  0, 38),
                ( 0, 34, 34, 34, 34, 34,  0, 38),
                (34, 34, 34, 34, 34, 34, 34, 38)
        )),
        (   handle => FOREST_TILE_BITMAP,
            bitmap => (
                (11, 11, 11, 11, 12,  1, 11, 11),
                (12,  1, 11, 11, 11, 12, 11, 11),
                (11, 12, 11, 11, 11, 11, 11, 11),
                (11, 11, 11, 12, 11, 11, 11, 11),
                (11, 11, 11, 11, 12, 11, 11, 11),
                (11, 11, 11, 11, 11, 11,  1, 11),
                (11, 12, 11, 11, 11, 11, 12, 11),
                (11, 11, 12, 11, 11, 11, 11, 11)
        )),
        (
            handle => GAME_OVER_TILE_BITMAP,
            bitmap => (
                (22, 46, 22, 46, 22, 46, 22, 22),
                (22, 22, 46, 26, 26, 26, 46, 22),
                (22, 46, 26, 53, 53, 53, 25, 22),
                (22, 26, 53, 53, 53, 53, 53, 42),
                (22, 42, 53, 53, 34, 53, 34, 23),
                (22, 22, 23, 36, 53, 34, 53, 23),
                (22, 22, 22, 23, 36, 36, 36, 23),
                (22, 22, 22, 22, 24, 23, 23, 22)
            )
        ),
        (
            handle => GAME_WON_TILE_BITMAP,
            bitmap => (
                ( 7,  7, 38, 38, 38, 38, 38,  7),
                ( 7,  7, 38, 46, 46,  1, 38, 17),
                ( 7,  7, 46, 26, 46, 46, 38, 17),
                ( 7, 46, 26, 46, 26, 46, 38,  7),
                (38, 38, 38, 38, 38, 38, 38,  7),
                (38,  1, 46,  2, 38,  2, 38,  7),
                (38,  2,  1,  2, 38,  2, 38,  7),
                (38, 38, 38, 38, 38, 38,  7,  7)
            )
        )
    );

end;
